library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use	IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity TEMPLATE is
	port (B : in STD_LOGIC;
		  A	: in STD_LOGIC;
		  Z : out STD_LOGIC);
end TEMPLATE;

architecture RTL of TEMPLATE is

begin

end RTL;