library ieee;
use ieee.std_logic_1164.all;
--use ieee.std_logic_arith.all;
--use ieee.std_logic_unsigned.all;

entity TEMPLATE is
	port ( A, B, C, D : in std_logic;
		   Z : out std_logic);
end TEMPLATE;

architecture Behavioral of TEMPLATE is

begin
	
end Behavioral;